module memory 
#(
    parameter A = 12,  // Address width
    parameter m = 16   // Data width
)
(
    input CLK,                   // Clock signal
    input [A-1:0] address,       // Memory address
    input [m-1:0] data_in,       // Data to write into memory
    input write_enable,          // Enable signal for write operation
    input read_enable,           // Enable signal for read operation
    output [m-1:0] data_out  // Data read from memory
);
    localparam D = (1 << A);  // Number of memory locations (2^A)
    reg [m-1:0] mem [0:D-1];  // Memory array

    // Initialize memory during simulation or provide default values
    initial begin
        // Initializing memory locations with non-zero values
        // memory initiailization for all machine codes used in the program 
		mem[16'h012c] = 16'h11f4;//Add
        mem[16'h012d] = 16'h01f5;//AND
        mem[16'h012e] = 16'h21f6;//LDA
        mem[16'h012f] = 16'h31f7;//STA
        mem[16'h0130] = 16'h4300;//BUN
        mem[16'h0131] = 16'h51f9;//BSA
        mem[16'h0132] = 16'h61fa;//ISZ
        mem[16'h0133] = 16'h81fb;//Add INDIRECT
        mem[16'h0134] = 16'h91fc;//AND INDIRECT
        mem[16'h0135] = 16'ha1fd;//LDA INDIRECT
        mem[16'h0136] = 16'hb1fe;//STA INDIRECT
        mem[16'h0137] = 16'hc1ff;//BUN INDIRECT
        mem[16'h0138] = 16'hd200;//BSA INDIRECT
        mem[16'h0139] = 16'he201;//ISZ INDIRECT
        mem[16'h013a] = 16'h7800;//CLA
        mem[16'h013b] = 16'h7400;//CLE
        mem[16'h013c] = 16'h7200;//CMA
        mem[16'h013d] = 16'h7100;//CME
        mem[16'h013e] = 16'h7080;//CIR
        mem[16'h013f] = 16'h7040;//CIL
        mem[16'h0140] = 16'h7020;//INC
        mem[16'h0141] = 16'h7010;//SPA
        mem[16'h0142] = 16'h7008;//SNA
        mem[16'h0143] = 16'h7004;//SZA
        mem[16'h0144] = 16'h7002;//SZE
        mem[16'h0145] = 16'h7001;//HLT
        //////////////////////////////
        //////////////////////////////
        mem[16'h0146] = 16'hf800;//INP
        mem[16'h0147] = 16'hf400;//OUT
        mem[16'h0148] = 16'hf200;//SKI
        mem[16'h0149] = 16'hf100;//SKO
        mem[16'h014a] = 16'hf080;//ION
        mem[16'h014b] = 16'hf040;//IOF
		// memory initialization for the values used in the DR for the memory reference instructions
        mem[16'h01f4] = 16'h1010;
        mem[16'h01f5] = 16'h0101;
        mem[16'h01f6] = 16'h1234;
        mem[16'h01f7] = 16'h0000;
        mem[16'h01f8] = 16'h014a;
        mem[16'h01f9] = 16'h014b;
        mem[16'h01fa] = 16'h4132;
        mem[16'h01fb] = 16'h0258;
        mem[16'h01fc] = 16'h0259;
        mem[16'h01fd] = 16'h025a;
        mem[16'h01fe] = 16'h025b;
        mem[16'h01ff] = 16'h025c;
        mem[16'h0200] = 16'h0400;
        mem[16'h0201] = 16'h025e;
		//memory initialization for the values used in the DR for the memory reference instructions
		mem[16'h0258] = 16'h1010;
        mem[16'h0259] = 16'h0101;
        mem[16'h025a] = 16'h1234;
        mem[16'h025b] = 16'h0000;
        mem[16'h025c] = 16'h4138;
        mem[16'h025d] = 16'h014B;
        mem[16'h025e] = 16'h0000;
        mem[16'h025f] = 16'h0000;
        mem[16'h0300] = 16'h4131;
	    mem[16'h0400] = 16'h4139;
		mem[16'h0401] = 16'h4139;
		

    end

    always @(posedge CLK) begin
        if (write_enable) begin
            mem[address] = data_in;  // Write data to the memory
        end

        
    end
	assign data_out = (read_enable)? mem[address]: 16'bx;

	
	
endmodule